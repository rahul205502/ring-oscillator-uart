`timescale 1ns/1ps

module edge_detector ( input clk, input ro_out,input rst_n, output edge_dec );

    reg ro_out_prev;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin 
            ro_out_prev <= 1'b0;
        end
        else begin 
            ro_out_prev <= ro_out ;
        end
     end
     
     assign edge_dec = (~ro_out_prev) & ro_out ;
endmodule